module ysyx_22041461_IF(
  input  wire [63:0] pc  ,
  output wire [31:0] inst
);